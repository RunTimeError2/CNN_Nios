// kernel.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module kernel (
		input  wire        clk_clk,                                         //                        clk.clk
		inout  wire [7:0]  lcd1602_demo_conduit_end_0_export_data,          // lcd1602_demo_conduit_end_0.export_data
		output wire        lcd1602_demo_conduit_end_0_export_rw,            //                           .export_rw
		output wire        lcd1602_demo_conduit_end_0_export_en,            //                           .export_en
		output wire        lcd1602_demo_conduit_end_0_export_rs,            //                           .export_rs
		output wire        lcd1602_demo_conduit_end_0_export_blon,          //                           .export_blon
		output wire        lcd1602_demo_conduit_end_0_export_on,            //                           .export_on
		output wire        pio_external_connection_export,                  //    pio_external_connection.export
		input  wire        reset_reset_n,                                   //                      reset.reset_n
		output wire [12:0] sdram_controller_wire_addr,                      //      sdram_controller_wire.addr
		output wire [1:0]  sdram_controller_wire_ba,                        //                           .ba
		output wire        sdram_controller_wire_cas_n,                     //                           .cas_n
		output wire        sdram_controller_wire_cke,                       //                           .cke
		output wire        sdram_controller_wire_cs_n,                      //                           .cs_n
		inout  wire [31:0] sdram_controller_wire_dq,                        //                           .dq
		output wire [3:0]  sdram_controller_wire_dqm,                       //                           .dqm
		output wire        sdram_controller_wire_ras_n,                     //                           .ras_n
		output wire        sdram_controller_wire_we_n,                      //                           .we_n
		output wire        user_gio_pwm_conduit_end_0_export,               // user_gio_pwm_conduit_end_0.export
		input  wire        user_ir_conduit_end_0_export_input,              //      user_ir_conduit_end_0.export_input
		input  wire        user_ltm_adc_conduit_end_0_export_irst_n,        // user_ltm_adc_conduit_end_0.export_irst_n
		output wire        user_ltm_adc_conduit_end_0_export_oadc_din,      //                           .export_oadc_din
		output wire        user_ltm_adc_conduit_end_0_export_oadc_dclk,     //                           .export_oadc_dclk
		output wire        user_ltm_adc_conduit_end_0_export_oadc_cs,       //                           .export_oadc_cs
		input  wire        user_ltm_adc_conduit_end_0_export_iadc_dout,     //                           .export_iadc_dout
		input  wire        user_ltm_adc_conduit_end_0_export_iadc_busy,     //                           .export_iadc_busy
		input  wire        user_ltm_adc_conduit_end_0_export_iadc_penirq_n, //                           .export_iadc_penirq_n
		output wire        user_ltm_adc_conduit_end_0_export_otouch_irq,    //                           .export_otouch_irq
		output wire [6:0]  user_seg8_conduit_end_0_export_0,                //    user_seg8_conduit_end_0.export_0
		output wire [6:0]  user_seg8_conduit_end_0_export_1,                //                           .export_1
		output wire [6:0]  user_seg8_conduit_end_0_export_2,                //                           .export_2
		output wire [6:0]  user_seg8_conduit_end_0_export_3,                //                           .export_3
		output wire [6:0]  user_seg8_conduit_end_0_export_4,                //                           .export_4
		output wire [6:0]  user_seg8_conduit_end_0_export_5,                //                           .export_5
		output wire [6:0]  user_seg8_conduit_end_0_export_6,                //                           .export_6
		output wire [6:0]  user_seg8_conduit_end_0_export_7,                //                           .export_7
		output wire [19:0] user_sram_bw_conduit_end_0_export_osram_addr,    // user_sram_bw_conduit_end_0.export_osram_addr
		inout  wire [15:0] user_sram_bw_conduit_end_0_export_iosram_dq,     //                           .export_iosram_dq
		output wire        user_sram_bw_conduit_end_0_export_osram_we_n,    //                           .export_osram_we_n
		output wire        user_sram_bw_conduit_end_0_export_osram_oe_n,    //                           .export_osram_oe_n
		output wire        user_sram_bw_conduit_end_0_export_osram_ub_n,    //                           .export_osram_ub_n
		output wire        user_sram_bw_conduit_end_0_export_osram_lb_n,    //                           .export_osram_lb_n
		output wire        user_sram_bw_conduit_end_0_export_osram_ce_n,    //                           .export_osram_ce_n
		input  wire        user_sram_bw_conduit_end_0_export_irst_n,        //                           .export_irst_n
		output wire [31:0] user_sram_bw_conduit_end_0_export_osram_data,    //                           .export_osram_data
		input  wire        user_sram_bw_conduit_end_0_export_iread_sram_en, //                           .export_iread_sram_en
		input  wire        user_sram_bw_conduit_end_0_export_iclk50m        //                           .export_iclk50m
	);

	wire  [31:0] nios2_data_master_readdata;                                // mm_interconnect_0:nios2_data_master_readdata -> nios2:d_readdata
	wire         nios2_data_master_waitrequest;                             // mm_interconnect_0:nios2_data_master_waitrequest -> nios2:d_waitrequest
	wire         nios2_data_master_debugaccess;                             // nios2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_data_master_debugaccess
	wire  [28:0] nios2_data_master_address;                                 // nios2:d_address -> mm_interconnect_0:nios2_data_master_address
	wire   [3:0] nios2_data_master_byteenable;                              // nios2:d_byteenable -> mm_interconnect_0:nios2_data_master_byteenable
	wire         nios2_data_master_read;                                    // nios2:d_read -> mm_interconnect_0:nios2_data_master_read
	wire         nios2_data_master_write;                                   // nios2:d_write -> mm_interconnect_0:nios2_data_master_write
	wire  [31:0] nios2_data_master_writedata;                               // nios2:d_writedata -> mm_interconnect_0:nios2_data_master_writedata
	wire  [31:0] nios2_instruction_master_readdata;                         // mm_interconnect_0:nios2_instruction_master_readdata -> nios2:i_readdata
	wire         nios2_instruction_master_waitrequest;                      // mm_interconnect_0:nios2_instruction_master_waitrequest -> nios2:i_waitrequest
	wire  [28:0] nios2_instruction_master_address;                          // nios2:i_address -> mm_interconnect_0:nios2_instruction_master_address
	wire         nios2_instruction_master_read;                             // nios2:i_read -> mm_interconnect_0:nios2_instruction_master_read
	wire         nios2_instruction_master_readdatavalid;                    // mm_interconnect_0:nios2_instruction_master_readdatavalid -> nios2:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_0_user_gio_pwm_avalon_slave_0_chipselect;  // mm_interconnect_0:User_GIO_PWM_avalon_slave_0_chipselect -> User_GIO_PWM:avs_chipselect
	wire  [31:0] mm_interconnect_0_user_gio_pwm_avalon_slave_0_readdata;    // User_GIO_PWM:avs_readdata -> mm_interconnect_0:User_GIO_PWM_avalon_slave_0_readdata
	wire   [3:0] mm_interconnect_0_user_gio_pwm_avalon_slave_0_address;     // mm_interconnect_0:User_GIO_PWM_avalon_slave_0_address -> User_GIO_PWM:avs_address
	wire         mm_interconnect_0_user_gio_pwm_avalon_slave_0_read;        // mm_interconnect_0:User_GIO_PWM_avalon_slave_0_read -> User_GIO_PWM:avs_read
	wire         mm_interconnect_0_user_gio_pwm_avalon_slave_0_write;       // mm_interconnect_0:User_GIO_PWM_avalon_slave_0_write -> User_GIO_PWM:avs_write
	wire  [31:0] mm_interconnect_0_user_gio_pwm_avalon_slave_0_writedata;   // mm_interconnect_0:User_GIO_PWM_avalon_slave_0_writedata -> User_GIO_PWM:avs_writedata
	wire         mm_interconnect_0_lcd1602_demo_avalon_slave_0_chipselect;  // mm_interconnect_0:LCD1602_Demo_avalon_slave_0_chipselect -> LCD1602_Demo:avs_chipselect
	wire  [31:0] mm_interconnect_0_lcd1602_demo_avalon_slave_0_readdata;    // LCD1602_Demo:avs_readdata -> mm_interconnect_0:LCD1602_Demo_avalon_slave_0_readdata
	wire   [4:0] mm_interconnect_0_lcd1602_demo_avalon_slave_0_address;     // mm_interconnect_0:LCD1602_Demo_avalon_slave_0_address -> LCD1602_Demo:avs_address
	wire         mm_interconnect_0_lcd1602_demo_avalon_slave_0_read;        // mm_interconnect_0:LCD1602_Demo_avalon_slave_0_read -> LCD1602_Demo:avs_read
	wire         mm_interconnect_0_lcd1602_demo_avalon_slave_0_write;       // mm_interconnect_0:LCD1602_Demo_avalon_slave_0_write -> LCD1602_Demo:avs_write
	wire  [31:0] mm_interconnect_0_lcd1602_demo_avalon_slave_0_writedata;   // mm_interconnect_0:LCD1602_Demo_avalon_slave_0_writedata -> LCD1602_Demo:avs_writedata
	wire         mm_interconnect_0_user_ir_avalon_slave_0_chipselect;       // mm_interconnect_0:User_IR_avalon_slave_0_chipselect -> User_IR:avs_chipselect
	wire  [31:0] mm_interconnect_0_user_ir_avalon_slave_0_readdata;         // User_IR:avs_readdata -> mm_interconnect_0:User_IR_avalon_slave_0_readdata
	wire   [3:0] mm_interconnect_0_user_ir_avalon_slave_0_address;          // mm_interconnect_0:User_IR_avalon_slave_0_address -> User_IR:avs_address
	wire         mm_interconnect_0_user_ir_avalon_slave_0_read;             // mm_interconnect_0:User_IR_avalon_slave_0_read -> User_IR:avs_read
	wire         mm_interconnect_0_user_ir_avalon_slave_0_write;            // mm_interconnect_0:User_IR_avalon_slave_0_write -> User_IR:avs_write
	wire  [31:0] mm_interconnect_0_user_ir_avalon_slave_0_writedata;        // mm_interconnect_0:User_IR_avalon_slave_0_writedata -> User_IR:avs_writedata
	wire         mm_interconnect_0_user_seg8_avalon_slave_0_chipselect;     // mm_interconnect_0:User_SEG8_avalon_slave_0_chipselect -> User_SEG8:avs_chipselect
	wire  [31:0] mm_interconnect_0_user_seg8_avalon_slave_0_readdata;       // User_SEG8:avs_readdata -> mm_interconnect_0:User_SEG8_avalon_slave_0_readdata
	wire   [3:0] mm_interconnect_0_user_seg8_avalon_slave_0_address;        // mm_interconnect_0:User_SEG8_avalon_slave_0_address -> User_SEG8:avs_address
	wire         mm_interconnect_0_user_seg8_avalon_slave_0_read;           // mm_interconnect_0:User_SEG8_avalon_slave_0_read -> User_SEG8:avs_read
	wire         mm_interconnect_0_user_seg8_avalon_slave_0_write;          // mm_interconnect_0:User_SEG8_avalon_slave_0_write -> User_SEG8:avs_write
	wire  [31:0] mm_interconnect_0_user_seg8_avalon_slave_0_writedata;      // mm_interconnect_0:User_SEG8_avalon_slave_0_writedata -> User_SEG8:avs_writedata
	wire         mm_interconnect_0_user_ltm_adc_avalon_slave_0_chipselect;  // mm_interconnect_0:User_LTM_ADC_avalon_slave_0_chipselect -> User_LTM_ADC:avs_chipselect
	wire  [31:0] mm_interconnect_0_user_ltm_adc_avalon_slave_0_readdata;    // User_LTM_ADC:avs_readdata -> mm_interconnect_0:User_LTM_ADC_avalon_slave_0_readdata
	wire   [3:0] mm_interconnect_0_user_ltm_adc_avalon_slave_0_address;     // mm_interconnect_0:User_LTM_ADC_avalon_slave_0_address -> User_LTM_ADC:avs_address
	wire         mm_interconnect_0_user_ltm_adc_avalon_slave_0_read;        // mm_interconnect_0:User_LTM_ADC_avalon_slave_0_read -> User_LTM_ADC:avs_read
	wire         mm_interconnect_0_user_ltm_adc_avalon_slave_0_write;       // mm_interconnect_0:User_LTM_ADC_avalon_slave_0_write -> User_LTM_ADC:avs_write
	wire  [31:0] mm_interconnect_0_user_ltm_adc_avalon_slave_0_writedata;   // mm_interconnect_0:User_LTM_ADC_avalon_slave_0_writedata -> User_LTM_ADC:avs_writedata
	wire         mm_interconnect_0_user_sram_bw_avalon_slave_0_chipselect;  // mm_interconnect_0:User_SRAM_BW_avalon_slave_0_chipselect -> User_SRAM_BW:avs_chipselect
	wire  [31:0] mm_interconnect_0_user_sram_bw_avalon_slave_0_readdata;    // User_SRAM_BW:avs_readdata -> mm_interconnect_0:User_SRAM_BW_avalon_slave_0_readdata
	wire   [3:0] mm_interconnect_0_user_sram_bw_avalon_slave_0_address;     // mm_interconnect_0:User_SRAM_BW_avalon_slave_0_address -> User_SRAM_BW:avs_address
	wire         mm_interconnect_0_user_sram_bw_avalon_slave_0_read;        // mm_interconnect_0:User_SRAM_BW_avalon_slave_0_read -> User_SRAM_BW:avs_read
	wire         mm_interconnect_0_user_sram_bw_avalon_slave_0_write;       // mm_interconnect_0:User_SRAM_BW_avalon_slave_0_write -> User_SRAM_BW:avs_write
	wire  [31:0] mm_interconnect_0_user_sram_bw_avalon_slave_0_writedata;   // mm_interconnect_0:User_SRAM_BW_avalon_slave_0_writedata -> User_SRAM_BW:avs_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;       // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;        // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_readdata;          // nios2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_debug_mem_slave_waitrequest;       // nios2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_debug_mem_slave_debugaccess;       // mm_interconnect_0:nios2_debug_mem_slave_debugaccess -> nios2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_debug_mem_slave_address;           // mm_interconnect_0:nios2_debug_mem_slave_address -> nios2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_debug_mem_slave_read;              // mm_interconnect_0:nios2_debug_mem_slave_read -> nios2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_debug_mem_slave_byteenable;        // mm_interconnect_0:nios2_debug_mem_slave_byteenable -> nios2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_debug_mem_slave_write;             // mm_interconnect_0:nios2_debug_mem_slave_write -> nios2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_writedata;         // mm_interconnect_0:nios2_debug_mem_slave_writedata -> nios2:debug_mem_slave_writedata
	wire         mm_interconnect_0_sdram_controller_s1_chipselect;          // mm_interconnect_0:sdram_controller_s1_chipselect -> sdram_controller:az_cs
	wire  [31:0] mm_interconnect_0_sdram_controller_s1_readdata;            // sdram_controller:za_data -> mm_interconnect_0:sdram_controller_s1_readdata
	wire         mm_interconnect_0_sdram_controller_s1_waitrequest;         // sdram_controller:za_waitrequest -> mm_interconnect_0:sdram_controller_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_controller_s1_address;             // mm_interconnect_0:sdram_controller_s1_address -> sdram_controller:az_addr
	wire         mm_interconnect_0_sdram_controller_s1_read;                // mm_interconnect_0:sdram_controller_s1_read -> sdram_controller:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_controller_s1_byteenable;          // mm_interconnect_0:sdram_controller_s1_byteenable -> sdram_controller:az_be_n
	wire         mm_interconnect_0_sdram_controller_s1_readdatavalid;       // sdram_controller:za_valid -> mm_interconnect_0:sdram_controller_s1_readdatavalid
	wire         mm_interconnect_0_sdram_controller_s1_write;               // mm_interconnect_0:sdram_controller_s1_write -> sdram_controller:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_controller_s1_writedata;           // mm_interconnect_0:sdram_controller_s1_writedata -> sdram_controller:az_data
	wire         mm_interconnect_0_pio_s1_chipselect;                       // mm_interconnect_0:pio_s1_chipselect -> pio:chipselect
	wire  [31:0] mm_interconnect_0_pio_s1_readdata;                         // pio:readdata -> mm_interconnect_0:pio_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_s1_address;                          // mm_interconnect_0:pio_s1_address -> pio:address
	wire         mm_interconnect_0_pio_s1_write;                            // mm_interconnect_0:pio_s1_write -> pio:write_n
	wire  [31:0] mm_interconnect_0_pio_s1_writedata;                        // mm_interconnect_0:pio_s1_writedata -> pio:writedata
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // User_IR:avs_irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_irq_irq;                                             // irq_mapper:sender_irq -> nios2:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [LCD1602_Demo:csi_RST_N, User_GIO_PWM:csi_reset_n, User_IR:csi_reset_n, User_LTM_ADC:csi_reset_n, User_SEG8:csi_reset_n, User_SRAM_BW:csi_reset_n, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:nios2_reset_reset_bridge_in_reset_reset, nios2:reset_n, pio:reset_n, rst_translator:in_reset, sdram_controller:reset_n, sysid_qsys:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [nios2:reset_req, rst_translator:reset_req_in]
	wire         nios2_debug_reset_request_reset;                           // nios2:debug_reset_request -> rst_controller:reset_in1

	LCD_Module lcd1602_demo (
		.csi_CLK        (clk_clk),                                                  //          clock.clk
		.csi_RST_N      (~rst_controller_reset_out_reset),                          //    clock_reset.reset_n
		.avs_chipselect (mm_interconnect_0_lcd1602_demo_avalon_slave_0_chipselect), // avalon_slave_0.chipselect
		.avs_address    (mm_interconnect_0_lcd1602_demo_avalon_slave_0_address),    //               .address
		.avs_read       (mm_interconnect_0_lcd1602_demo_avalon_slave_0_read),       //               .read
		.avs_readdata   (mm_interconnect_0_lcd1602_demo_avalon_slave_0_readdata),   //               .readdata
		.avs_write      (mm_interconnect_0_lcd1602_demo_avalon_slave_0_write),      //               .write
		.avs_writedata  (mm_interconnect_0_lcd1602_demo_avalon_slave_0_writedata),  //               .writedata
		.coe_LCD_DATA   (lcd1602_demo_conduit_end_0_export_data),                   //  conduit_end_0.export_data
		.coe_LCD_RW     (lcd1602_demo_conduit_end_0_export_rw),                     //               .export_rw
		.coe_LCD_EN     (lcd1602_demo_conduit_end_0_export_en),                     //               .export_en
		.coe_LCD_RS     (lcd1602_demo_conduit_end_0_export_rs),                     //               .export_rs
		.coe_LCD_BLON   (lcd1602_demo_conduit_end_0_export_blon),                   //               .export_blon
		.coe_LCD_ON     (lcd1602_demo_conduit_end_0_export_on)                      //               .export_on
	);

	User_Demo user_gio_pwm (
		.avs_chipselect (mm_interconnect_0_user_gio_pwm_avalon_slave_0_chipselect), // avalon_slave_0.chipselect
		.avs_address    (mm_interconnect_0_user_gio_pwm_avalon_slave_0_address),    //               .address
		.avs_read       (mm_interconnect_0_user_gio_pwm_avalon_slave_0_read),       //               .read
		.avs_readdata   (mm_interconnect_0_user_gio_pwm_avalon_slave_0_readdata),   //               .readdata
		.avs_write      (mm_interconnect_0_user_gio_pwm_avalon_slave_0_write),      //               .write
		.avs_writedata  (mm_interconnect_0_user_gio_pwm_avalon_slave_0_writedata),  //               .writedata
		.csi_clk        (clk_clk),                                                  //          clock.clk
		.csi_reset_n    (~rst_controller_reset_out_reset),                          //    clock_reset.reset_n
		.coe_GPIO_LED   (user_gio_pwm_conduit_end_0_export)                         //  conduit_end_0.export
	);

	IR_Module #(
		.IDLE              (3'b000),
		.GUIDANCE          (3'b001),
		.DATAREAD          (3'b010),
		.IDLE_HIGH_DUR     (262143),
		.GUIDE_LOW_DUR     (230000),
		.GUIDE_HIGH_DUR    (210000),
		.DATA_HIGH_DUR     (41500),
		.BIT_AVAILABLE_DUR (20000)
	) user_ir (
		.csi_clk          (clk_clk),                                             //          clock.clk
		.csi_reset_n      (~rst_controller_reset_out_reset),                     //    clock_reset.reset_n
		.avs_chipselect   (mm_interconnect_0_user_ir_avalon_slave_0_chipselect), // avalon_slave_0.chipselect
		.avs_address      (mm_interconnect_0_user_ir_avalon_slave_0_address),    //               .address
		.avs_read         (mm_interconnect_0_user_ir_avalon_slave_0_read),       //               .read
		.avs_readdata     (mm_interconnect_0_user_ir_avalon_slave_0_readdata),   //               .readdata
		.avs_write        (mm_interconnect_0_user_ir_avalon_slave_0_write),      //               .write
		.avs_writedata    (mm_interconnect_0_user_ir_avalon_slave_0_writedata),  //               .writedata
		.avs_irq          (irq_mapper_receiver1_irq),                            //            irq.irq
		.coe_IRData_Input (user_ir_conduit_end_0_export_input)                   //  conduit_end_0.export_input
	);

	adc_spi_controller #(
		.SYSCLK_FRQ   (50000000),
		.ADC_DCLK_FRQ (1000)
	) user_ltm_adc (
		.csi_clk           (clk_clk),                                                  //          clock.clk
		.csi_reset_n       (~rst_controller_reset_out_reset),                          //    clock_reset.reset_n
		.avs_chipselect    (mm_interconnect_0_user_ltm_adc_avalon_slave_0_chipselect), // avalon_slave_0.chipselect
		.avs_address       (mm_interconnect_0_user_ltm_adc_avalon_slave_0_address),    //               .address
		.avs_read          (mm_interconnect_0_user_ltm_adc_avalon_slave_0_read),       //               .read
		.avs_readdata      (mm_interconnect_0_user_ltm_adc_avalon_slave_0_readdata),   //               .readdata
		.avs_write         (mm_interconnect_0_user_ltm_adc_avalon_slave_0_write),      //               .write
		.avs_writedata     (mm_interconnect_0_user_ltm_adc_avalon_slave_0_writedata),  //               .writedata
		.coe_iRST_n        (user_ltm_adc_conduit_end_0_export_irst_n),                 //  conduit_end_0.export_irst_n
		.coe_oADC_DIN      (user_ltm_adc_conduit_end_0_export_oadc_din),               //               .export_oadc_din
		.coe_oADC_DCLK     (user_ltm_adc_conduit_end_0_export_oadc_dclk),              //               .export_oadc_dclk
		.coe_oADC_CS       (user_ltm_adc_conduit_end_0_export_oadc_cs),                //               .export_oadc_cs
		.coe_iADC_DOUT     (user_ltm_adc_conduit_end_0_export_iadc_dout),              //               .export_iadc_dout
		.coe_iADC_BUSY     (user_ltm_adc_conduit_end_0_export_iadc_busy),              //               .export_iadc_busy
		.coe_iADC_PENIRQ_n (user_ltm_adc_conduit_end_0_export_iadc_penirq_n),          //               .export_iadc_penirq_n
		.coe_oTOUCH_IRQ    (user_ltm_adc_conduit_end_0_export_otouch_irq)              //               .export_otouch_irq
	);

	SEG7_LUT_8 user_seg8 (
		.csi_clk        (clk_clk),                                               //          clock.clk
		.csi_reset_n    (~rst_controller_reset_out_reset),                       //    clock_reset.reset_n
		.avs_chipselect (mm_interconnect_0_user_seg8_avalon_slave_0_chipselect), // avalon_slave_0.chipselect
		.avs_address    (mm_interconnect_0_user_seg8_avalon_slave_0_address),    //               .address
		.avs_read       (mm_interconnect_0_user_seg8_avalon_slave_0_read),       //               .read
		.avs_readdata   (mm_interconnect_0_user_seg8_avalon_slave_0_readdata),   //               .readdata
		.avs_write      (mm_interconnect_0_user_seg8_avalon_slave_0_write),      //               .write
		.avs_writedata  (mm_interconnect_0_user_seg8_avalon_slave_0_writedata),  //               .writedata
		.coe_oSEG0      (user_seg8_conduit_end_0_export_0),                      //  conduit_end_0.export_0
		.coe_oSEG1      (user_seg8_conduit_end_0_export_1),                      //               .export_1
		.coe_oSEG2      (user_seg8_conduit_end_0_export_2),                      //               .export_2
		.coe_oSEG3      (user_seg8_conduit_end_0_export_3),                      //               .export_3
		.coe_oSEG4      (user_seg8_conduit_end_0_export_4),                      //               .export_4
		.coe_oSEG5      (user_seg8_conduit_end_0_export_5),                      //               .export_5
		.coe_oSEG6      (user_seg8_conduit_end_0_export_6),                      //               .export_6
		.coe_oSEG7      (user_seg8_conduit_end_0_export_7)                       //               .export_7
	);

	SRAM_Image_BW user_sram_bw (
		.csi_clk           (clk_clk),                                                  //          clock.clk
		.csi_reset_n       (~rst_controller_reset_out_reset),                          //    clock_reset.reset_n
		.avs_chipselect    (mm_interconnect_0_user_sram_bw_avalon_slave_0_chipselect), // avalon_slave_0.chipselect
		.avs_address       (mm_interconnect_0_user_sram_bw_avalon_slave_0_address),    //               .address
		.avs_read          (mm_interconnect_0_user_sram_bw_avalon_slave_0_read),       //               .read
		.avs_readdata      (mm_interconnect_0_user_sram_bw_avalon_slave_0_readdata),   //               .readdata
		.avs_write         (mm_interconnect_0_user_sram_bw_avalon_slave_0_write),      //               .write
		.avs_writedata     (mm_interconnect_0_user_sram_bw_avalon_slave_0_writedata),  //               .writedata
		.coe_oSRAM_ADDR    (user_sram_bw_conduit_end_0_export_osram_addr),             //  conduit_end_0.export_osram_addr
		.coe_ioSRAM_DQ     (user_sram_bw_conduit_end_0_export_iosram_dq),              //               .export_iosram_dq
		.coe_oSRAM_WE_N    (user_sram_bw_conduit_end_0_export_osram_we_n),             //               .export_osram_we_n
		.coe_oSRAM_OE_N    (user_sram_bw_conduit_end_0_export_osram_oe_n),             //               .export_osram_oe_n
		.coe_oSRAM_UB_N    (user_sram_bw_conduit_end_0_export_osram_ub_n),             //               .export_osram_ub_n
		.coe_oSRAM_LB_N    (user_sram_bw_conduit_end_0_export_osram_lb_n),             //               .export_osram_lb_n
		.coe_oSRAM_CE_N    (user_sram_bw_conduit_end_0_export_osram_ce_n),             //               .export_osram_ce_n
		.coe_iRST_n        (user_sram_bw_conduit_end_0_export_irst_n),                 //               .export_irst_n
		.coe_oSRAM_DATA    (user_sram_bw_conduit_end_0_export_osram_data),             //               .export_osram_data
		.coe_iREAD_SRAM_EN (user_sram_bw_conduit_end_0_export_iread_sram_en),          //               .export_iread_sram_en
		.coe_iCLK50M       (user_sram_bw_conduit_end_0_export_iclk50m)                 //               .export_iclk50m
	);

	kernel_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	kernel_nios2 nios2 (
		.clk                                 (clk_clk),                                             //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (nios2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                     // custom_instruction_master.readra
	);

	kernel_pio pio (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_s1_readdata),   //                    .readdata
		.out_port   (pio_external_connection_export)       // external_connection.export
	);

	kernel_sdram_controller sdram_controller (
		.clk            (clk_clk),                                             //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                     // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_controller_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_controller_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_controller_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_controller_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_controller_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_controller_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_controller_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_controller_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_controller_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_controller_wire_addr),                          //  wire.export
		.zs_ba          (sdram_controller_wire_ba),                            //      .export
		.zs_cas_n       (sdram_controller_wire_cas_n),                         //      .export
		.zs_cke         (sdram_controller_wire_cke),                           //      .export
		.zs_cs_n        (sdram_controller_wire_cs_n),                          //      .export
		.zs_dq          (sdram_controller_wire_dq),                            //      .export
		.zs_dqm         (sdram_controller_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_controller_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_controller_wire_we_n)                           //      .export
	);

	kernel_sysid_qsys sysid_qsys (
		.clock    (clk_clk),                                             //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	kernel_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                             (clk_clk),                                                   //                           clk_clk.clk
		.nios2_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // nios2_reset_reset_bridge_in_reset.reset
		.nios2_data_master_address               (nios2_data_master_address),                                 //                 nios2_data_master.address
		.nios2_data_master_waitrequest           (nios2_data_master_waitrequest),                             //                                  .waitrequest
		.nios2_data_master_byteenable            (nios2_data_master_byteenable),                              //                                  .byteenable
		.nios2_data_master_read                  (nios2_data_master_read),                                    //                                  .read
		.nios2_data_master_readdata              (nios2_data_master_readdata),                                //                                  .readdata
		.nios2_data_master_write                 (nios2_data_master_write),                                   //                                  .write
		.nios2_data_master_writedata             (nios2_data_master_writedata),                               //                                  .writedata
		.nios2_data_master_debugaccess           (nios2_data_master_debugaccess),                             //                                  .debugaccess
		.nios2_instruction_master_address        (nios2_instruction_master_address),                          //          nios2_instruction_master.address
		.nios2_instruction_master_waitrequest    (nios2_instruction_master_waitrequest),                      //                                  .waitrequest
		.nios2_instruction_master_read           (nios2_instruction_master_read),                             //                                  .read
		.nios2_instruction_master_readdata       (nios2_instruction_master_readdata),                         //                                  .readdata
		.nios2_instruction_master_readdatavalid  (nios2_instruction_master_readdatavalid),                    //                                  .readdatavalid
		.jtag_uart_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //       jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                  .write
		.jtag_uart_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                  .read
		.jtag_uart_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                  .readdata
		.jtag_uart_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                  .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                  .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                  .chipselect
		.LCD1602_Demo_avalon_slave_0_address     (mm_interconnect_0_lcd1602_demo_avalon_slave_0_address),     //       LCD1602_Demo_avalon_slave_0.address
		.LCD1602_Demo_avalon_slave_0_write       (mm_interconnect_0_lcd1602_demo_avalon_slave_0_write),       //                                  .write
		.LCD1602_Demo_avalon_slave_0_read        (mm_interconnect_0_lcd1602_demo_avalon_slave_0_read),        //                                  .read
		.LCD1602_Demo_avalon_slave_0_readdata    (mm_interconnect_0_lcd1602_demo_avalon_slave_0_readdata),    //                                  .readdata
		.LCD1602_Demo_avalon_slave_0_writedata   (mm_interconnect_0_lcd1602_demo_avalon_slave_0_writedata),   //                                  .writedata
		.LCD1602_Demo_avalon_slave_0_chipselect  (mm_interconnect_0_lcd1602_demo_avalon_slave_0_chipselect),  //                                  .chipselect
		.nios2_debug_mem_slave_address           (mm_interconnect_0_nios2_debug_mem_slave_address),           //             nios2_debug_mem_slave.address
		.nios2_debug_mem_slave_write             (mm_interconnect_0_nios2_debug_mem_slave_write),             //                                  .write
		.nios2_debug_mem_slave_read              (mm_interconnect_0_nios2_debug_mem_slave_read),              //                                  .read
		.nios2_debug_mem_slave_readdata          (mm_interconnect_0_nios2_debug_mem_slave_readdata),          //                                  .readdata
		.nios2_debug_mem_slave_writedata         (mm_interconnect_0_nios2_debug_mem_slave_writedata),         //                                  .writedata
		.nios2_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_debug_mem_slave_byteenable),        //                                  .byteenable
		.nios2_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_debug_mem_slave_waitrequest),       //                                  .waitrequest
		.nios2_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_debug_mem_slave_debugaccess),       //                                  .debugaccess
		.pio_s1_address                          (mm_interconnect_0_pio_s1_address),                          //                            pio_s1.address
		.pio_s1_write                            (mm_interconnect_0_pio_s1_write),                            //                                  .write
		.pio_s1_readdata                         (mm_interconnect_0_pio_s1_readdata),                         //                                  .readdata
		.pio_s1_writedata                        (mm_interconnect_0_pio_s1_writedata),                        //                                  .writedata
		.pio_s1_chipselect                       (mm_interconnect_0_pio_s1_chipselect),                       //                                  .chipselect
		.sdram_controller_s1_address             (mm_interconnect_0_sdram_controller_s1_address),             //               sdram_controller_s1.address
		.sdram_controller_s1_write               (mm_interconnect_0_sdram_controller_s1_write),               //                                  .write
		.sdram_controller_s1_read                (mm_interconnect_0_sdram_controller_s1_read),                //                                  .read
		.sdram_controller_s1_readdata            (mm_interconnect_0_sdram_controller_s1_readdata),            //                                  .readdata
		.sdram_controller_s1_writedata           (mm_interconnect_0_sdram_controller_s1_writedata),           //                                  .writedata
		.sdram_controller_s1_byteenable          (mm_interconnect_0_sdram_controller_s1_byteenable),          //                                  .byteenable
		.sdram_controller_s1_readdatavalid       (mm_interconnect_0_sdram_controller_s1_readdatavalid),       //                                  .readdatavalid
		.sdram_controller_s1_waitrequest         (mm_interconnect_0_sdram_controller_s1_waitrequest),         //                                  .waitrequest
		.sdram_controller_s1_chipselect          (mm_interconnect_0_sdram_controller_s1_chipselect),          //                                  .chipselect
		.sysid_qsys_control_slave_address        (mm_interconnect_0_sysid_qsys_control_slave_address),        //          sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata       (mm_interconnect_0_sysid_qsys_control_slave_readdata),       //                                  .readdata
		.User_GIO_PWM_avalon_slave_0_address     (mm_interconnect_0_user_gio_pwm_avalon_slave_0_address),     //       User_GIO_PWM_avalon_slave_0.address
		.User_GIO_PWM_avalon_slave_0_write       (mm_interconnect_0_user_gio_pwm_avalon_slave_0_write),       //                                  .write
		.User_GIO_PWM_avalon_slave_0_read        (mm_interconnect_0_user_gio_pwm_avalon_slave_0_read),        //                                  .read
		.User_GIO_PWM_avalon_slave_0_readdata    (mm_interconnect_0_user_gio_pwm_avalon_slave_0_readdata),    //                                  .readdata
		.User_GIO_PWM_avalon_slave_0_writedata   (mm_interconnect_0_user_gio_pwm_avalon_slave_0_writedata),   //                                  .writedata
		.User_GIO_PWM_avalon_slave_0_chipselect  (mm_interconnect_0_user_gio_pwm_avalon_slave_0_chipselect),  //                                  .chipselect
		.User_IR_avalon_slave_0_address          (mm_interconnect_0_user_ir_avalon_slave_0_address),          //            User_IR_avalon_slave_0.address
		.User_IR_avalon_slave_0_write            (mm_interconnect_0_user_ir_avalon_slave_0_write),            //                                  .write
		.User_IR_avalon_slave_0_read             (mm_interconnect_0_user_ir_avalon_slave_0_read),             //                                  .read
		.User_IR_avalon_slave_0_readdata         (mm_interconnect_0_user_ir_avalon_slave_0_readdata),         //                                  .readdata
		.User_IR_avalon_slave_0_writedata        (mm_interconnect_0_user_ir_avalon_slave_0_writedata),        //                                  .writedata
		.User_IR_avalon_slave_0_chipselect       (mm_interconnect_0_user_ir_avalon_slave_0_chipselect),       //                                  .chipselect
		.User_LTM_ADC_avalon_slave_0_address     (mm_interconnect_0_user_ltm_adc_avalon_slave_0_address),     //       User_LTM_ADC_avalon_slave_0.address
		.User_LTM_ADC_avalon_slave_0_write       (mm_interconnect_0_user_ltm_adc_avalon_slave_0_write),       //                                  .write
		.User_LTM_ADC_avalon_slave_0_read        (mm_interconnect_0_user_ltm_adc_avalon_slave_0_read),        //                                  .read
		.User_LTM_ADC_avalon_slave_0_readdata    (mm_interconnect_0_user_ltm_adc_avalon_slave_0_readdata),    //                                  .readdata
		.User_LTM_ADC_avalon_slave_0_writedata   (mm_interconnect_0_user_ltm_adc_avalon_slave_0_writedata),   //                                  .writedata
		.User_LTM_ADC_avalon_slave_0_chipselect  (mm_interconnect_0_user_ltm_adc_avalon_slave_0_chipselect),  //                                  .chipselect
		.User_SEG8_avalon_slave_0_address        (mm_interconnect_0_user_seg8_avalon_slave_0_address),        //          User_SEG8_avalon_slave_0.address
		.User_SEG8_avalon_slave_0_write          (mm_interconnect_0_user_seg8_avalon_slave_0_write),          //                                  .write
		.User_SEG8_avalon_slave_0_read           (mm_interconnect_0_user_seg8_avalon_slave_0_read),           //                                  .read
		.User_SEG8_avalon_slave_0_readdata       (mm_interconnect_0_user_seg8_avalon_slave_0_readdata),       //                                  .readdata
		.User_SEG8_avalon_slave_0_writedata      (mm_interconnect_0_user_seg8_avalon_slave_0_writedata),      //                                  .writedata
		.User_SEG8_avalon_slave_0_chipselect     (mm_interconnect_0_user_seg8_avalon_slave_0_chipselect),     //                                  .chipselect
		.User_SRAM_BW_avalon_slave_0_address     (mm_interconnect_0_user_sram_bw_avalon_slave_0_address),     //       User_SRAM_BW_avalon_slave_0.address
		.User_SRAM_BW_avalon_slave_0_write       (mm_interconnect_0_user_sram_bw_avalon_slave_0_write),       //                                  .write
		.User_SRAM_BW_avalon_slave_0_read        (mm_interconnect_0_user_sram_bw_avalon_slave_0_read),        //                                  .read
		.User_SRAM_BW_avalon_slave_0_readdata    (mm_interconnect_0_user_sram_bw_avalon_slave_0_readdata),    //                                  .readdata
		.User_SRAM_BW_avalon_slave_0_writedata   (mm_interconnect_0_user_sram_bw_avalon_slave_0_writedata),   //                                  .writedata
		.User_SRAM_BW_avalon_slave_0_chipselect  (mm_interconnect_0_user_sram_bw_avalon_slave_0_chipselect)   //                                  .chipselect
	);

	kernel_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios2_debug_reset_request_reset),    // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
